package util is
	TYPE andar IS (andar0, andar1, andar2, andar3, andar4, andar5, andar6);
end util;